`define BIAS_FILE_0_0 "mifs/b_0_0.mif"
`define WEIGHT_FILE_0_0 "mifs/w_0_0.mif"
`define BIAS_FILE_0_1 "mifs/b_0_1.mif"
`define WEIGHT_FILE_0_1 "mifs/w_0_1.mif"
`define BIAS_FILE_0_2 "mifs/b_0_2.mif"
`define WEIGHT_FILE_0_2 "mifs/w_0_2.mif"
`define BIAS_FILE_0_3 "mifs/b_0_3.mif"
`define WEIGHT_FILE_0_3 "mifs/w_0_3.mif"
`define BIAS_FILE_0_4 "mifs/b_0_4.mif"
`define WEIGHT_FILE_0_4 "mifs/w_0_4.mif"
`define BIAS_FILE_0_5 "mifs/b_0_5.mif"
`define WEIGHT_FILE_0_5 "mifs/w_0_5.mif"
`define BIAS_FILE_0_6 "mifs/b_0_6.mif"
`define WEIGHT_FILE_0_6 "mifs/w_0_6.mif"
`define BIAS_FILE_0_7 "mifs/b_0_7.mif"
`define WEIGHT_FILE_0_7 "mifs/w_0_7.mif"
`define BIAS_FILE_0_8 "mifs/b_0_8.mif"
`define WEIGHT_FILE_0_8 "mifs/w_0_8.mif"
`define BIAS_FILE_0_9 "mifs/b_0_9.mif"
`define WEIGHT_FILE_0_9 "mifs/w_0_9.mif"
`define BIAS_FILE_0_10 "mifs/b_0_10.mif"
`define WEIGHT_FILE_0_10 "mifs/w_0_10.mif"
`define BIAS_FILE_0_11 "mifs/b_0_11.mif"
`define WEIGHT_FILE_0_11 "mifs/w_0_11.mif"
`define BIAS_FILE_0_12 "mifs/b_0_12.mif"
`define WEIGHT_FILE_0_12 "mifs/w_0_12.mif"
`define BIAS_FILE_0_13 "mifs/b_0_13.mif"
`define WEIGHT_FILE_0_13 "mifs/w_0_13.mif"
`define BIAS_FILE_0_14 "mifs/b_0_14.mif"
`define WEIGHT_FILE_0_14 "mifs/w_0_14.mif"
`define BIAS_FILE_0_15 "mifs/b_0_15.mif"
`define WEIGHT_FILE_0_15 "mifs/w_0_15.mif"
`define BIAS_FILE_0_16 "mifs/b_0_16.mif"
`define WEIGHT_FILE_0_16 "mifs/w_0_16.mif"
`define BIAS_FILE_0_17 "mifs/b_0_17.mif"
`define WEIGHT_FILE_0_17 "mifs/w_0_17.mif"
`define BIAS_FILE_0_18 "mifs/b_0_18.mif"
`define WEIGHT_FILE_0_18 "mifs/w_0_18.mif"
`define BIAS_FILE_0_19 "mifs/b_0_19.mif"
`define WEIGHT_FILE_0_19 "mifs/w_0_19.mif"
`define BIAS_FILE_0_20 "mifs/b_0_20.mif"
`define WEIGHT_FILE_0_20 "mifs/w_0_20.mif"
`define BIAS_FILE_0_21 "mifs/b_0_21.mif"
`define WEIGHT_FILE_0_21 "mifs/w_0_21.mif"
`define BIAS_FILE_0_22 "mifs/b_0_22.mif"
`define WEIGHT_FILE_0_22 "mifs/w_0_22.mif"
`define BIAS_FILE_0_23 "mifs/b_0_23.mif"
`define WEIGHT_FILE_0_23 "mifs/w_0_23.mif"
`define BIAS_FILE_0_24 "mifs/b_0_24.mif"
`define WEIGHT_FILE_0_24 "mifs/w_0_24.mif"
`define BIAS_FILE_0_25 "mifs/b_0_25.mif"
`define WEIGHT_FILE_0_25 "mifs/w_0_25.mif"
`define BIAS_FILE_0_26 "mifs/b_0_26.mif"
`define WEIGHT_FILE_0_26 "mifs/w_0_26.mif"
`define BIAS_FILE_0_27 "mifs/b_0_27.mif"
`define WEIGHT_FILE_0_27 "mifs/w_0_27.mif"
`define BIAS_FILE_0_28 "mifs/b_0_28.mif"
`define WEIGHT_FILE_0_28 "mifs/w_0_28.mif"
`define BIAS_FILE_0_29 "mifs/b_0_29.mif"
`define WEIGHT_FILE_0_29 "mifs/w_0_29.mif"
`define BIAS_FILE_1_0 "mifs/b_1_0.mif"
`define WEIGHT_FILE_1_0 "mifs/w_1_0.mif"
`define BIAS_FILE_1_1 "mifs/b_1_1.mif"
`define WEIGHT_FILE_1_1 "mifs/w_1_1.mif"
`define BIAS_FILE_1_2 "mifs/b_1_2.mif"
`define WEIGHT_FILE_1_2 "mifs/w_1_2.mif"
`define BIAS_FILE_1_3 "mifs/b_1_3.mif"
`define WEIGHT_FILE_1_3 "mifs/w_1_3.mif"
`define BIAS_FILE_1_4 "mifs/b_1_4.mif"
`define WEIGHT_FILE_1_4 "mifs/w_1_4.mif"
`define BIAS_FILE_1_5 "mifs/b_1_5.mif"
`define WEIGHT_FILE_1_5 "mifs/w_1_5.mif"
`define BIAS_FILE_1_6 "mifs/b_1_6.mif"
`define WEIGHT_FILE_1_6 "mifs/w_1_6.mif"
`define BIAS_FILE_1_7 "mifs/b_1_7.mif"
`define WEIGHT_FILE_1_7 "mifs/w_1_7.mif"
`define BIAS_FILE_1_8 "mifs/b_1_8.mif"
`define WEIGHT_FILE_1_8 "mifs/w_1_8.mif"
`define BIAS_FILE_1_9 "mifs/b_1_9.mif"
`define WEIGHT_FILE_1_9 "mifs/w_1_9.mif"
`define BIAS_FILE_1_10 "mifs/b_1_10.mif"
`define WEIGHT_FILE_1_10 "mifs/w_1_10.mif"
`define BIAS_FILE_1_11 "mifs/b_1_11.mif"
`define WEIGHT_FILE_1_11 "mifs/w_1_11.mif"
`define BIAS_FILE_1_12 "mifs/b_1_12.mif"
`define WEIGHT_FILE_1_12 "mifs/w_1_12.mif"
`define BIAS_FILE_1_13 "mifs/b_1_13.mif"
`define WEIGHT_FILE_1_13 "mifs/w_1_13.mif"
`define BIAS_FILE_1_14 "mifs/b_1_14.mif"
`define WEIGHT_FILE_1_14 "mifs/w_1_14.mif"
`define BIAS_FILE_1_15 "mifs/b_1_15.mif"
`define WEIGHT_FILE_1_15 "mifs/w_1_15.mif"
`define BIAS_FILE_1_16 "mifs/b_1_16.mif"
`define WEIGHT_FILE_1_16 "mifs/w_1_16.mif"
`define BIAS_FILE_1_17 "mifs/b_1_17.mif"
`define WEIGHT_FILE_1_17 "mifs/w_1_17.mif"
`define BIAS_FILE_1_18 "mifs/b_1_18.mif"
`define WEIGHT_FILE_1_18 "mifs/w_1_18.mif"
`define BIAS_FILE_1_19 "mifs/b_1_19.mif"
`define WEIGHT_FILE_1_19 "mifs/w_1_19.mif"
`define BIAS_FILE_1_20 "mifs/b_1_20.mif"
`define WEIGHT_FILE_1_20 "mifs/w_1_20.mif"
`define BIAS_FILE_1_21 "mifs/b_1_21.mif"
`define WEIGHT_FILE_1_21 "mifs/w_1_21.mif"
`define BIAS_FILE_1_22 "mifs/b_1_22.mif"
`define WEIGHT_FILE_1_22 "mifs/w_1_22.mif"
`define BIAS_FILE_1_23 "mifs/b_1_23.mif"
`define WEIGHT_FILE_1_23 "mifs/w_1_23.mif"
`define BIAS_FILE_1_24 "mifs/b_1_24.mif"
`define WEIGHT_FILE_1_24 "mifs/w_1_24.mif"
`define BIAS_FILE_1_25 "mifs/b_1_25.mif"
`define WEIGHT_FILE_1_25 "mifs/w_1_25.mif"
`define BIAS_FILE_1_26 "mifs/b_1_26.mif"
`define WEIGHT_FILE_1_26 "mifs/w_1_26.mif"
`define BIAS_FILE_1_27 "mifs/b_1_27.mif"
`define WEIGHT_FILE_1_27 "mifs/w_1_27.mif"
`define BIAS_FILE_1_28 "mifs/b_1_28.mif"
`define WEIGHT_FILE_1_28 "mifs/w_1_28.mif"
`define BIAS_FILE_1_29 "mifs/b_1_29.mif"
`define WEIGHT_FILE_1_29 "mifs/w_1_29.mif"
`define BIAS_FILE_2_0 "mifs/b_2_0.mif"
`define WEIGHT_FILE_2_0 "mifs/w_2_0.mif"
`define BIAS_FILE_2_1 "mifs/b_2_1.mif"
`define WEIGHT_FILE_2_1 "mifs/w_2_1.mif"
`define BIAS_FILE_2_2 "mifs/b_2_2.mif"
`define WEIGHT_FILE_2_2 "mifs/w_2_2.mif"
`define BIAS_FILE_2_3 "mifs/b_2_3.mif"
`define WEIGHT_FILE_2_3 "mifs/w_2_3.mif"
`define BIAS_FILE_2_4 "mifs/b_2_4.mif"
`define WEIGHT_FILE_2_4 "mifs/w_2_4.mif"
`define BIAS_FILE_2_5 "mifs/b_2_5.mif"
`define WEIGHT_FILE_2_5 "mifs/w_2_5.mif"
`define BIAS_FILE_2_6 "mifs/b_2_6.mif"
`define WEIGHT_FILE_2_6 "mifs/w_2_6.mif"
`define BIAS_FILE_2_7 "mifs/b_2_7.mif"
`define WEIGHT_FILE_2_7 "mifs/w_2_7.mif"
`define BIAS_FILE_2_8 "mifs/b_2_8.mif"
`define WEIGHT_FILE_2_8 "mifs/w_2_8.mif"
`define BIAS_FILE_2_9 "mifs/b_2_9.mif"
`define WEIGHT_FILE_2_9 "mifs/w_2_9.mif"
`define BIAS_FILE_3_0 "mifs/b_3_0.mif"
`define WEIGHT_FILE_3_0 "mifs/w_3_0.mif"
