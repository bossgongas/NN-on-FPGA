`define BIAS_FILE_0_0 "b_0_0.mif"
`define WEIGHT_FILE_0_0 "w_0_0.mif"
`define BIAS_FILE_0_1 "b_0_1.mif"
`define WEIGHT_FILE_0_1 "w_0_1.mif"
`define BIAS_FILE_0_2 "b_0_2.mif"
`define WEIGHT_FILE_0_2 "w_0_2.mif"
`define BIAS_FILE_0_3 "b_0_3.mif"
`define WEIGHT_FILE_0_3 "w_0_3.mif"
`define BIAS_FILE_0_4 "b_0_4.mif"
`define WEIGHT_FILE_0_4 "w_0_4.mif"
`define BIAS_FILE_0_5 "b_0_5.mif"
`define WEIGHT_FILE_0_5 "w_0_5.mif"
`define BIAS_FILE_0_6 "b_0_6.mif"
`define WEIGHT_FILE_0_6 "w_0_6.mif"
`define BIAS_FILE_0_7 "b_0_7.mif"
`define WEIGHT_FILE_0_7 "w_0_7.mif"
`define BIAS_FILE_0_8 "b_0_8.mif"
`define WEIGHT_FILE_0_8 "w_0_8.mif"
`define BIAS_FILE_0_9 "b_0_9.mif"
`define WEIGHT_FILE_0_9 "w_0_9.mif"
`define BIAS_FILE_0_10 "b_0_10.mif"
`define WEIGHT_FILE_0_10 "w_0_10.mif"
`define BIAS_FILE_0_11 "b_0_11.mif"
`define WEIGHT_FILE_0_11 "w_0_11.mif"
`define BIAS_FILE_0_12 "b_0_12.mif"
`define WEIGHT_FILE_0_12 "w_0_12.mif"
`define BIAS_FILE_0_13 "b_0_13.mif"
`define WEIGHT_FILE_0_13 "w_0_13.mif"
`define BIAS_FILE_0_14 "b_0_14.mif"
`define WEIGHT_FILE_0_14 "w_0_14.mif"
`define BIAS_FILE_0_15 "b_0_15.mif"
`define WEIGHT_FILE_0_15 "w_0_15.mif"
`define BIAS_FILE_0_16 "b_0_16.mif"
`define WEIGHT_FILE_0_16 "w_0_16.mif"
`define BIAS_FILE_0_17 "b_0_17.mif"
`define WEIGHT_FILE_0_17 "w_0_17.mif"
`define BIAS_FILE_0_18 "b_0_18.mif"
`define WEIGHT_FILE_0_18 "w_0_18.mif"
`define BIAS_FILE_0_19 "b_0_19.mif"
`define WEIGHT_FILE_0_19 "w_0_19.mif"
`define BIAS_FILE_0_20 "b_0_20.mif"
`define WEIGHT_FILE_0_20 "w_0_20.mif"
`define BIAS_FILE_0_21 "b_0_21.mif"
`define WEIGHT_FILE_0_21 "w_0_21.mif"
`define BIAS_FILE_0_22 "b_0_22.mif"
`define WEIGHT_FILE_0_22 "w_0_22.mif"
`define BIAS_FILE_0_23 "b_0_23.mif"
`define WEIGHT_FILE_0_23 "w_0_23.mif"
`define BIAS_FILE_0_24 "b_0_24.mif"
`define WEIGHT_FILE_0_24 "w_0_24.mif"
`define BIAS_FILE_0_25 "b_0_25.mif"
`define WEIGHT_FILE_0_25 "w_0_25.mif"
`define BIAS_FILE_0_26 "b_0_26.mif"
`define WEIGHT_FILE_0_26 "w_0_26.mif"
`define BIAS_FILE_0_27 "b_0_27.mif"
`define WEIGHT_FILE_0_27 "w_0_27.mif"
`define BIAS_FILE_0_28 "b_0_28.mif"
`define WEIGHT_FILE_0_28 "w_0_28.mif"
`define BIAS_FILE_0_29 "b_0_29.mif"
`define WEIGHT_FILE_0_29 "w_0_29.mif"
`define BIAS_FILE_1_0 "b_1_0.mif"
`define WEIGHT_FILE_1_0 "w_1_0.mif"
`define BIAS_FILE_1_1 "b_1_1.mif"
`define WEIGHT_FILE_1_1 "w_1_1.mif"
`define BIAS_FILE_1_2 "b_1_2.mif"
`define WEIGHT_FILE_1_2 "w_1_2.mif"
`define BIAS_FILE_1_3 "b_1_3.mif"
`define WEIGHT_FILE_1_3 "w_1_3.mif"
`define BIAS_FILE_1_4 "b_1_4.mif"
`define WEIGHT_FILE_1_4 "w_1_4.mif"
`define BIAS_FILE_1_5 "b_1_5.mif"
`define WEIGHT_FILE_1_5 "w_1_5.mif"
`define BIAS_FILE_1_6 "b_1_6.mif"
`define WEIGHT_FILE_1_6 "w_1_6.mif"
`define BIAS_FILE_1_7 "b_1_7.mif"
`define WEIGHT_FILE_1_7 "w_1_7.mif"
`define BIAS_FILE_1_8 "b_1_8.mif"
`define WEIGHT_FILE_1_8 "w_1_8.mif"
`define BIAS_FILE_1_9 "b_1_9.mif"
`define WEIGHT_FILE_1_9 "w_1_9.mif"
`define BIAS_FILE_1_10 "b_1_10.mif"
`define WEIGHT_FILE_1_10 "w_1_10.mif"
`define BIAS_FILE_1_11 "b_1_11.mif"
`define WEIGHT_FILE_1_11 "w_1_11.mif"
`define BIAS_FILE_1_12 "b_1_12.mif"
`define WEIGHT_FILE_1_12 "w_1_12.mif"
`define BIAS_FILE_1_13 "b_1_13.mif"
`define WEIGHT_FILE_1_13 "w_1_13.mif"
`define BIAS_FILE_1_14 "b_1_14.mif"
`define WEIGHT_FILE_1_14 "w_1_14.mif"
`define BIAS_FILE_1_15 "b_1_15.mif"
`define WEIGHT_FILE_1_15 "w_1_15.mif"
`define BIAS_FILE_1_16 "b_1_16.mif"
`define WEIGHT_FILE_1_16 "w_1_16.mif"
`define BIAS_FILE_1_17 "b_1_17.mif"
`define WEIGHT_FILE_1_17 "w_1_17.mif"
`define BIAS_FILE_1_18 "b_1_18.mif"
`define WEIGHT_FILE_1_18 "w_1_18.mif"
`define BIAS_FILE_1_19 "b_1_19.mif"
`define WEIGHT_FILE_1_19 "w_1_19.mif"
`define BIAS_FILE_1_20 "b_1_20.mif"
`define WEIGHT_FILE_1_20 "w_1_20.mif"
`define BIAS_FILE_1_21 "b_1_21.mif"
`define WEIGHT_FILE_1_21 "w_1_21.mif"
`define BIAS_FILE_1_22 "b_1_22.mif"
`define WEIGHT_FILE_1_22 "w_1_22.mif"
`define BIAS_FILE_1_23 "b_1_23.mif"
`define WEIGHT_FILE_1_23 "w_1_23.mif"
`define BIAS_FILE_1_24 "b_1_24.mif"
`define WEIGHT_FILE_1_24 "w_1_24.mif"
`define BIAS_FILE_1_25 "b_1_25.mif"
`define WEIGHT_FILE_1_25 "w_1_25.mif"
`define BIAS_FILE_1_26 "b_1_26.mif"
`define WEIGHT_FILE_1_26 "w_1_26.mif"
`define BIAS_FILE_1_27 "b_1_27.mif"
`define WEIGHT_FILE_1_27 "w_1_27.mif"
`define BIAS_FILE_1_28 "b_1_28.mif"
`define WEIGHT_FILE_1_28 "w_1_28.mif"
`define BIAS_FILE_1_29 "b_1_29.mif"
`define WEIGHT_FILE_1_29 "w_1_29.mif"
`define BIAS_FILE_2_0 "b_2_0.mif"
`define WEIGHT_FILE_2_0 "w_2_0.mif"
`define BIAS_FILE_2_1 "b_2_1.mif"
`define WEIGHT_FILE_2_1 "w_2_1.mif"
`define BIAS_FILE_2_2 "b_2_2.mif"
`define WEIGHT_FILE_2_2 "w_2_2.mif"
`define BIAS_FILE_2_3 "b_2_3.mif"
`define WEIGHT_FILE_2_3 "w_2_3.mif"
`define BIAS_FILE_2_4 "b_2_4.mif"
`define WEIGHT_FILE_2_4 "w_2_4.mif"
`define BIAS_FILE_2_5 "b_2_5.mif"
`define WEIGHT_FILE_2_5 "w_2_5.mif"
`define BIAS_FILE_2_6 "b_2_6.mif"
`define WEIGHT_FILE_2_6 "w_2_6.mif"
`define BIAS_FILE_2_7 "b_2_7.mif"
`define WEIGHT_FILE_2_7 "w_2_7.mif"
`define BIAS_FILE_2_8 "b_2_8.mif"
`define WEIGHT_FILE_2_8 "w_2_8.mif"
`define BIAS_FILE_2_9 "b_2_9.mif"
`define WEIGHT_FILE_2_9 "w_2_9.mif"
`define BIAS_FILE_3_0 "b_3_0.mif"
`define WEIGHT_FILE_3_0 "w_3_0.mif"
